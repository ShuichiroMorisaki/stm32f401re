
signature sADC {
};

celltype tADC {
	entry sADC eADC;
};